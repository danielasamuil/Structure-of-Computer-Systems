----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/12/2020 07:29:14 PM
-- Design Name: 
-- Module Name: CarryBlock - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CarryBlock is
generic (n: integer);
port (x: in std_logic_vector (n downto 0);
y: in std_logic_vector (n downto 0);
C0: in std_logic;
C: out std_logic );
end CarryBlock;

architecture Behavioral of CarryBlock is 

signal aux_carry1: std_logic;
signal aux_carry2: std_logic;
signal aux_carry3: std_logic;
signal aux_carry4: std_logic;
signal aux_carry5: std_logic;
signal aux_carry6: std_logic;
signal aux_carry7: std_logic;
signal aux_carry8: std_logic;
signal aux_carry9: std_logic;
signal aux_carry10: std_logic;
signal aux_carry11: std_logic;
signal aux_carry12: std_logic;
signal aux_carry13: std_logic;
signal aux_carry14: std_logic;
signal aux_carry15: std_logic;

begin

process (x,y,C0)
begin

if (n=0) then 
C <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
elsif (n=1) then 
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
C <= (x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1));
elsif (n=2) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
C <= (x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2));
elsif (n=3) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
C <= (x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3));
elsif (n=4) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
C <= (x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4));
elsif (n=5) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
C <= (x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5));
elsif (n=6) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
C <= (x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6));
elsif (n=7) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
C <= (x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7));
elsif (n=8) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
C <= (x(8) AND y(8)) OR (((x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7))) AND x(8)) OR (((x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7))) AND y(8));
elsif (n=9) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
C <= (x(9) AND y(9)) OR (((x(8) AND y(8)) OR (((x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7))) AND x(8)) OR (((x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7))) AND y(8))) AND x(9)) OR (((x(8) AND y(8)) OR (((x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7))) AND x(8)) OR (((x(7) AND y(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND x(7)) OR (((x(6) AND y(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND x(6)) OR (((x(5) AND y(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND x(5)) OR (((x(4) AND y(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND x(4)) OR (((x(3) AND y(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND x(3)) OR (((x(2) AND y(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND x(2)) OR (((x(1) AND y(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND x(1)) OR (((x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0))) AND y(1))) AND y(2))) AND y(3))) AND y(4))) AND y(5))) AND y(6))) AND y(7))) AND y(8))) AND y(9));
elsif (n=10) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
aux_carry10 <= (x(9) AND y(9)) OR (aux_carry9 AND x(9)) OR (aux_carry9 AND y(9));
C <= (x(10) AND y(10)) OR (x(10) AND aux_carry10) OR (y(10) AND aux_carry10);
elsif (n=11) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
aux_carry10 <= (x(9) AND y(9)) OR (aux_carry9 AND x(9)) OR (aux_carry9 AND y(9));
aux_carry11 <= (x(10) AND y(10)) OR (aux_carry10 AND x(10)) OR (aux_carry10 AND y(10));
C <= (x(11) AND y(11)) OR (aux_carry11 AND x(11)) OR (aux_carry11 AND y(11));
elsif (n=12) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND y(0)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
aux_carry10 <= (x(9) AND y(9)) OR (aux_carry9 AND x(9)) OR (aux_carry9 AND y(9));
aux_carry11 <= (x(10) AND y(10)) OR (aux_carry10 AND x(10)) OR (aux_carry10 AND y(10));
aux_carry12 <= (x(11) AND y(11)) OR (aux_carry11 AND x(11)) OR (aux_carry11 AND y(11));
C <= (x(12) AND y(12)) OR (aux_carry12 AND x(12)) OR (aux_carry12 AND y(12));
elsif (n=13) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
aux_carry10 <= (x(9) AND y(9)) OR (aux_carry9 AND x(9)) OR (aux_carry9 AND y(9));
aux_carry11 <= (x(10) AND y(10)) OR (aux_carry10 AND x(10)) OR (aux_carry10 AND y(10));
aux_carry12 <= (x(11) AND y(11)) OR (aux_carry11 AND x(11)) OR (aux_carry11 AND y(11));
aux_carry13 <= (x(12) AND y(12)) OR (aux_carry12 AND x(12)) OR (aux_carry12 AND y(12));
C <= (x(13) AND y(13)) OR (aux_carry13 AND x(13)) OR (aux_carry13 AND y(13));
elsif (n=14) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
aux_carry10 <= (x(9) AND y(9)) OR (aux_carry9 AND x(9)) OR (aux_carry9 AND y(9));
aux_carry11 <= (x(10) AND y(10)) OR (aux_carry10 AND x(10)) OR (aux_carry10 AND y(10));
aux_carry12 <= (x(11) AND y(11)) OR (aux_carry11 AND x(11)) OR (aux_carry11 AND y(11));
aux_carry13 <= (x(12) AND y(12)) OR (aux_carry12 AND x(12)) OR (aux_carry12 AND y(12));
aux_carry14 <= (x(13) AND y(13)) OR (aux_carry13 AND x(13)) OR (aux_carry13 AND y(13));
C <= (x(14) AND y(14)) OR (aux_carry14 AND x(14)) OR (aux_carry14 AND y(14));
elsif (n=15) then
aux_carry1 <= (x(0) AND y(0)) OR (C0 AND x(0)) OR (C0 AND y(0));
aux_carry2 <= (x(1) AND y(1)) OR (aux_carry1 AND x(1)) OR (aux_carry1 AND y(1));
aux_carry3 <= (x(2) AND y(2)) OR (aux_carry2 AND x(2)) OR (aux_carry2 AND y(2));
aux_carry4 <= (x(3) AND y(3)) OR (aux_carry3 AND x(3)) OR (aux_carry3 AND y(3));
aux_carry5 <= (x(4) AND y(4)) OR (aux_carry4 AND x(4)) OR (aux_carry4 AND y(4));
aux_carry6 <= (x(5) AND y(5)) OR (aux_carry5 AND x(5)) OR (aux_carry5 AND y(5));
aux_carry7 <= (x(6) AND y(6)) OR (aux_carry6 AND x(6)) OR (aux_carry6 AND y(6));
aux_carry8 <= (x(7) AND y(7)) OR (aux_carry7 AND x(7)) OR (aux_carry7 AND y(7));
aux_carry9 <= (x(8) AND y(8)) OR (aux_carry8 AND x(8)) OR (aux_carry8 AND y(8));
aux_carry10 <= (x(9) AND y(9)) OR (aux_carry9 AND x(9)) OR (aux_carry9 AND y(9));
aux_carry11 <= (x(10) AND y(10)) OR (aux_carry10 AND x(10)) OR (aux_carry10 AND y(10));
aux_carry12 <= (x(11) AND y(11)) OR (aux_carry11 AND x(11)) OR (aux_carry11 AND y(11));
aux_carry13 <= (x(12) AND y(12)) OR (aux_carry12 AND x(12)) OR (aux_carry12 AND y(12));
aux_carry14 <= (x(13) AND y(13)) OR (aux_carry13 AND x(13)) OR (aux_carry13 AND y(13));
aux_carry15 <= (x(14) AND y(14)) OR (aux_carry14 AND x(14)) OR (aux_carry14 AND y(14));
C <= (x(15) AND y(15)) OR (x(15) AND aux_carry15) OR (y(15) AND aux_carry15);
end if;

end process;
end Behavioral;
