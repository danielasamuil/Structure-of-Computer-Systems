----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/13/2020 12:21:11 PM
-- Design Name: 
-- Module Name: MULTIPLY_component - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_signed.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity WallaceTree is
Port (A: in std_logic_vector(15 downto 0);
B: in std_logic_vector(15 downto 0);
O: out std_logic_vector(29 downto 0) );
end WallaceTree;

architecture Behavioral of WallaceTree is

component Full_Adder is
port(nr1,nr2: in std_logic;
CIN: in std_logic;
adder_out: out std_logic;
COUT: out std_logic);
end component;

signal P0_0: std_logic;
signal P0_1: std_logic;
signal P0_2: std_logic;
signal P0_3: std_logic;
signal P0_4: std_logic;
signal P0_5: std_logic;
signal P0_6: std_logic;
signal P0_7: std_logic;
signal P0_8: std_logic;
signal P0_9: std_logic;
signal P0_10: std_logic;
signal P0_11: std_logic;
signal P0_12: std_logic;
signal P0_13: std_logic;
signal P0_14: std_logic;
signal P1_0: std_logic;
signal P1_1: std_logic;
signal P1_2: std_logic;
signal P1_3: std_logic;
signal P1_4: std_logic;
signal P1_5: std_logic;
signal P1_6: std_logic;
signal P1_7: std_logic;
signal P1_8: std_logic;
signal P1_9: std_logic;
signal P1_10: std_logic;
signal P1_11: std_logic;
signal P1_12: std_logic;
signal P1_13: std_logic;
signal P1_14: std_logic;
signal P2_0: std_logic;
signal P2_1: std_logic;
signal P2_2: std_logic;
signal P2_3: std_logic;
signal P2_4: std_logic;
signal P2_5: std_logic;
signal P2_6: std_logic;
signal P2_7: std_logic;
signal P2_8: std_logic;
signal P2_9: std_logic;
signal P2_10: std_logic;
signal P2_11: std_logic;
signal P2_12: std_logic;
signal P2_13: std_logic;
signal P2_14: std_logic;
signal P3_0: std_logic;
signal P3_1: std_logic;
signal P3_2: std_logic;
signal P3_3: std_logic;
signal P3_4: std_logic;
signal P3_5: std_logic;
signal P3_6: std_logic;
signal P3_7: std_logic;
signal P3_8: std_logic;
signal P3_9: std_logic;
signal P3_10: std_logic;
signal P3_11: std_logic;
signal P3_12: std_logic;
signal P3_13: std_logic;
signal P3_14: std_logic;
signal P4_0: std_logic;
signal P4_1: std_logic;
signal P4_2: std_logic;
signal P4_3: std_logic;
signal P4_4: std_logic;
signal P4_5: std_logic;
signal P4_6: std_logic;
signal P4_7: std_logic;
signal P4_8: std_logic;
signal P4_9: std_logic;
signal P4_10: std_logic;
signal P4_11: std_logic;
signal P4_12: std_logic;
signal P4_13: std_logic;
signal P4_14: std_logic;
signal P5_0: std_logic;
signal P5_1: std_logic;
signal P5_2: std_logic;
signal P5_3: std_logic;
signal P5_4: std_logic;
signal P5_5: std_logic;
signal P5_6: std_logic;
signal P5_7: std_logic;
signal P5_8: std_logic;
signal P5_9: std_logic;
signal P5_10: std_logic;
signal P5_11: std_logic;
signal P5_12: std_logic;
signal P5_13: std_logic;
signal P5_14: std_logic;
signal P6_0: std_logic;
signal P6_1: std_logic;
signal P6_2: std_logic;
signal P6_3: std_logic;
signal P6_4: std_logic;
signal P6_5: std_logic;
signal P6_6: std_logic;
signal P6_7: std_logic;
signal P6_8: std_logic;
signal P6_9: std_logic;
signal P6_10: std_logic;
signal P6_11: std_logic;
signal P6_12: std_logic;
signal P6_13: std_logic;
signal P6_14: std_logic;
signal P7_0: std_logic;
signal P7_1: std_logic;
signal P7_2: std_logic;
signal P7_3: std_logic;
signal P7_4: std_logic;
signal P7_5: std_logic;
signal P7_6: std_logic;
signal P7_7: std_logic;
signal P7_8: std_logic;
signal P7_9: std_logic;
signal P7_10: std_logic;
signal P7_11: std_logic;
signal P7_12: std_logic;
signal P7_13: std_logic;
signal P7_14: std_logic;
signal P8_0: std_logic;
signal P8_1: std_logic;
signal P8_2: std_logic;
signal P8_3: std_logic;
signal P8_4: std_logic;
signal P8_5: std_logic;
signal P8_6: std_logic;
signal P8_7: std_logic;
signal P8_8: std_logic;
signal P8_9: std_logic;
signal P8_10: std_logic;
signal P8_11: std_logic;
signal P8_12: std_logic;
signal P8_13: std_logic;
signal P8_14: std_logic;
signal P9_0: std_logic;
signal P9_1: std_logic;
signal P9_2: std_logic;
signal P9_3: std_logic;
signal P9_4: std_logic;
signal P9_5: std_logic;
signal P9_6: std_logic;
signal P9_7: std_logic;
signal P9_8: std_logic;
signal P9_9: std_logic;
signal P9_10: std_logic;
signal P9_11: std_logic;
signal P9_12: std_logic;
signal P9_13: std_logic;
signal P9_14: std_logic;
signal P10_0: std_logic;
signal P10_1: std_logic;
signal P10_2: std_logic;
signal P10_3: std_logic;
signal P10_4: std_logic;
signal P10_5: std_logic;
signal P10_6: std_logic;
signal P10_7: std_logic;
signal P10_8: std_logic;
signal P10_9: std_logic;
signal P10_10: std_logic;
signal P10_11: std_logic;
signal P10_12: std_logic;
signal P10_13: std_logic;
signal P10_14: std_logic;
signal P11_0: std_logic;
signal P11_1: std_logic;
signal P11_2: std_logic;
signal P11_3: std_logic;
signal P11_4: std_logic;
signal P11_5: std_logic;
signal P11_6: std_logic;
signal P11_7: std_logic;
signal P11_8: std_logic;
signal P11_9: std_logic;
signal P11_10: std_logic;
signal P11_11: std_logic;
signal P11_12: std_logic;
signal P11_13: std_logic;
signal P11_14: std_logic;
signal P12_0: std_logic;
signal P12_1: std_logic;
signal P12_2: std_logic;
signal P12_3: std_logic;
signal P12_4: std_logic;
signal P12_5: std_logic;
signal P12_6: std_logic;
signal P12_7: std_logic;
signal P12_8: std_logic;
signal P12_9: std_logic;
signal P12_10: std_logic;
signal P12_11: std_logic;
signal P12_12: std_logic;
signal P12_13: std_logic;
signal P12_14: std_logic;
signal P13_0: std_logic;
signal P13_1: std_logic;
signal P13_2: std_logic;
signal P13_3: std_logic;
signal P13_4: std_logic;
signal P13_5: std_logic;
signal P13_6: std_logic;
signal P13_7: std_logic;
signal P13_8: std_logic;
signal P13_9: std_logic;
signal P13_10: std_logic;
signal P13_11: std_logic;
signal P13_12: std_logic;
signal P13_13: std_logic;
signal P13_14: std_logic;
signal P14_0: std_logic;
signal P14_1: std_logic;
signal P14_2: std_logic;
signal P14_3: std_logic;
signal P14_4: std_logic;
signal P14_5: std_logic;
signal P14_6: std_logic;
signal P14_7: std_logic;
signal P14_8: std_logic;
signal P14_9: std_logic;
signal P14_10: std_logic;
signal P14_11: std_logic;
signal P14_12: std_logic;
signal P14_13: std_logic;
signal P14_14: std_logic;

signal C0: std_logic;
signal S0: std_logic;
signal C1: std_logic;
signal S1: std_logic;
signal C2: std_logic;
signal S2: std_logic;
signal C3: std_logic;
signal S3: std_logic;
signal C4: std_logic;
signal S4: std_logic;
signal C5: std_logic;
signal S5: std_logic;
signal C6: std_logic;
signal S6: std_logic;
signal C7: std_logic;
signal S7: std_logic;
signal C8: std_logic;
signal S8: std_logic;
signal C9: std_logic;
signal S9: std_logic;
signal C10: std_logic;
signal S10: std_logic;
signal C11: std_logic;
signal S11: std_logic;
signal C12: std_logic;
signal S12: std_logic;
signal C13: std_logic;
signal S13: std_logic;
signal C14: std_logic;
signal S14: std_logic;
signal C15: std_logic;
signal S15: std_logic;
signal C16: std_logic;
signal S16: std_logic;
signal C17: std_logic;
signal S17: std_logic;
signal C18: std_logic;
signal S18: std_logic;
signal C19: std_logic;
signal S19: std_logic;
signal C20: std_logic;
signal S20: std_logic;
signal C21: std_logic;
signal S21: std_logic;
signal C22: std_logic;
signal S22: std_logic;
signal C23: std_logic;
signal S23: std_logic;
signal C24: std_logic;
signal S24: std_logic;
signal C25: std_logic;
signal S25: std_logic;
signal C26: std_logic;
signal S26: std_logic;
signal C27: std_logic;
signal S27: std_logic;
signal C28: std_logic;
signal S28: std_logic;
signal C29: std_logic;
signal S29: std_logic;
signal C30: std_logic;
signal S30: std_logic;
signal C31: std_logic;
signal S31: std_logic;
signal C32: std_logic;
signal S32: std_logic;
signal C33: std_logic;
signal S33: std_logic;
signal C34: std_logic;
signal S34: std_logic;
signal C35: std_logic;
signal S35: std_logic;
signal C36: std_logic;
signal S36: std_logic;
signal C37: std_logic;
signal S37: std_logic;
signal C38: std_logic;
signal S38: std_logic;
signal C39: std_logic;
signal S39: std_logic;
signal C40: std_logic;
signal S40: std_logic;
signal C41: std_logic;
signal S41: std_logic;
signal C42: std_logic;
signal S42: std_logic;
signal C43: std_logic;
signal S43: std_logic;
signal C44: std_logic;
signal S44: std_logic;
signal C45: std_logic;
signal S45: std_logic;
signal C46: std_logic;
signal S46: std_logic;
signal C47: std_logic;
signal S47: std_logic;
signal C48: std_logic;
signal S48: std_logic;
signal C49: std_logic;
signal S49: std_logic;
signal C50: std_logic;
signal S50: std_logic;
signal C51: std_logic;
signal S51: std_logic;
signal C52: std_logic;
signal S52: std_logic;
signal C53: std_logic;
signal S53: std_logic;
signal C54: std_logic;
signal S54: std_logic;
signal C55: std_logic;
signal S55: std_logic;
signal C56: std_logic;
signal S56: std_logic;
signal C57: std_logic;
signal S57: std_logic;
signal C58: std_logic;
signal S58: std_logic;
signal C59: std_logic;
signal S59: std_logic;
signal C60: std_logic;
signal S60: std_logic;
signal C61: std_logic;
signal S61: std_logic;
signal C62: std_logic;
signal S62: std_logic;
signal C63: std_logic;
signal S63: std_logic;
signal C64: std_logic;
signal S64: std_logic;
signal C65: std_logic;
signal S65: std_logic;
signal C66: std_logic;
signal S66: std_logic;
signal C67: std_logic;
signal S67: std_logic;
signal C68: std_logic;
signal S68: std_logic;
signal C69: std_logic;
signal S69: std_logic;
signal C70: std_logic;
signal S70: std_logic;
signal C71: std_logic;
signal S71: std_logic;
signal C72: std_logic;
signal S72: std_logic;
signal C73: std_logic;
signal S73: std_logic;
signal C74: std_logic;
signal S74: std_logic;
signal C75: std_logic;
signal S75: std_logic;
signal C76: std_logic;
signal S76: std_logic;
signal C77: std_logic;
signal S77: std_logic;
signal C78: std_logic;
signal S78: std_logic;
signal C79: std_logic;
signal S79: std_logic;
signal C80: std_logic;
signal S80: std_logic;
signal C81: std_logic;
signal S81: std_logic;
signal C82: std_logic;
signal S82: std_logic;
signal C83: std_logic;
signal S83: std_logic;
signal C84: std_logic;
signal S84: std_logic;
signal C85: std_logic;
signal S85: std_logic;
signal C86: std_logic;
signal S86: std_logic;
signal C87: std_logic;
signal S87: std_logic;
signal C88: std_logic;
signal S88: std_logic;
signal C89: std_logic;
signal S89: std_logic;
signal C90: std_logic;
signal S90: std_logic;
signal C91: std_logic;
signal S91: std_logic;
signal C92: std_logic;
signal S92: std_logic;
signal C93: std_logic;
signal S93: std_logic;
signal C94: std_logic;
signal S94: std_logic;
signal C95: std_logic;
signal S95: std_logic;
signal C96: std_logic;
signal S96: std_logic;
signal C97: std_logic;
signal S97: std_logic;
signal C98: std_logic;
signal S98: std_logic;
signal C99: std_logic;
signal S99: std_logic;
signal C100: std_logic;
signal S100: std_logic;
signal C101: std_logic;
signal S101: std_logic;
signal C102: std_logic;
signal S102: std_logic;
signal C103: std_logic;
signal S103: std_logic;
signal C104: std_logic;
signal S104: std_logic;
signal C105: std_logic;
signal S105: std_logic;
signal C106: std_logic;
signal S106: std_logic;
signal C107: std_logic;
signal S107: std_logic;
signal C108: std_logic;
signal S108: std_logic;
signal C109: std_logic;
signal S109: std_logic;
signal C110: std_logic;
signal S110: std_logic;
signal C111: std_logic;
signal S111: std_logic;
signal C112: std_logic;
signal S112: std_logic;
signal C113: std_logic;
signal S113: std_logic;
signal C114: std_logic;
signal S114: std_logic;
signal C115: std_logic;
signal S115: std_logic;
signal C116: std_logic;
signal S116: std_logic;
signal C117: std_logic;
signal S117: std_logic;
signal C118: std_logic;
signal S118: std_logic;
signal C119: std_logic;
signal S119: std_logic;
signal C120: std_logic;
signal S120: std_logic;
signal C121: std_logic;
signal S121: std_logic;
signal C122: std_logic;
signal S122: std_logic;
signal C123: std_logic;
signal S123: std_logic;
signal C124: std_logic;
signal S124: std_logic;
signal C125: std_logic;
signal S125: std_logic;
signal C126: std_logic;
signal S126: std_logic;
signal C127: std_logic;
signal S127: std_logic;
signal C128: std_logic;
signal S128: std_logic;
signal C129: std_logic;
signal S129: std_logic;
signal C130: std_logic;
signal S130: std_logic;
signal C131: std_logic;
signal S131: std_logic;
signal C132: std_logic;
signal S132: std_logic;
signal C133: std_logic;
signal S133: std_logic;
signal C134: std_logic;
signal S134: std_logic;
signal C135: std_logic;
signal S135: std_logic;
signal C136: std_logic;
signal S136: std_logic;
signal C137: std_logic;
signal S137: std_logic;
signal C138: std_logic;
signal S138: std_logic;
signal C139: std_logic;
signal S139: std_logic;
signal C140: std_logic;
signal S140: std_logic;
signal C141: std_logic;
signal S141: std_logic;
signal C142: std_logic;
signal S142: std_logic;
signal C143: std_logic;
signal S143: std_logic;
signal C144: std_logic;
signal S144: std_logic;
signal C145: std_logic;
signal S145: std_logic;
signal C146: std_logic;
signal S146: std_logic;
signal C147: std_logic;
signal S147: std_logic;
signal C148: std_logic;
signal S148: std_logic;
signal C149: std_logic;
signal S149: std_logic;
signal C150: std_logic;
signal S150: std_logic;
signal C151: std_logic;
signal S151: std_logic;
signal C152: std_logic;
signal S152: std_logic;
signal C153: std_logic;
signal S153: std_logic;
signal C154: std_logic;
signal S154: std_logic;
signal C155: std_logic;
signal S155: std_logic;
signal C156: std_logic;
signal S156: std_logic;
signal C157: std_logic;
signal S157: std_logic;
signal C158: std_logic;
signal S158: std_logic;
signal C159: std_logic;
signal S159: std_logic;
signal C160: std_logic;
signal S160: std_logic;
signal C161: std_logic;
signal S161: std_logic;
signal C162: std_logic;
signal S162: std_logic;
signal C163: std_logic;
signal S163: std_logic;
signal C164: std_logic;
signal S164: std_logic;
signal C165: std_logic;
signal S165: std_logic;
signal C166: std_logic;
signal S166: std_logic;
signal C167: std_logic;
signal S167: std_logic;
signal C168: std_logic;
signal S168: std_logic;
signal C169: std_logic;
signal S169: std_logic;
signal C170: std_logic;
signal S170: std_logic;
signal C171: std_logic;
signal S171: std_logic;
signal C172: std_logic;
signal S172: std_logic;
signal C173: std_logic;
signal S173: std_logic;
signal C174: std_logic;
signal S174: std_logic;
signal C175: std_logic;
signal S175: std_logic;
signal C176: std_logic;
signal S176: std_logic;
signal C177: std_logic;
signal S177: std_logic;
signal C178: std_logic;
signal S178: std_logic;
signal C179: std_logic;
signal S179: std_logic;
signal C180: std_logic;
signal S180: std_logic;
signal C181: std_logic;
signal S181: std_logic;
signal C182: std_logic;
signal S182: std_logic;
signal C183: std_logic;
signal S183: std_logic;
signal C184: std_logic;
signal S184: std_logic;
signal C185: std_logic;
signal S185: std_logic;
signal C186: std_logic;
signal S186: std_logic;
signal C187: std_logic;
signal S187: std_logic;
signal C188: std_logic;
signal S188: std_logic;
signal C189: std_logic;
signal S189: std_logic;
signal C190: std_logic;
signal S190: std_logic;
signal C191: std_logic;
signal S191: std_logic;
signal C192: std_logic;
signal S192: std_logic;
signal C193: std_logic;
signal S193: std_logic;
signal C194: std_logic;
signal S194: std_logic;
signal C195: std_logic;
signal S195: std_logic;
signal C196: std_logic;
signal S196: std_logic;
signal C197: std_logic;
signal S197: std_logic;
signal C198: std_logic;
signal S198: std_logic;
signal C199: std_logic;
signal S199: std_logic;
signal C200: std_logic;
signal S200: std_logic;
signal C201: std_logic;
signal S201: std_logic;
signal C202: std_logic;
signal S202: std_logic;
signal C203: std_logic;
signal S203: std_logic;
signal C204: std_logic;
signal S204: std_logic;
signal C205: std_logic;
signal S205: std_logic;
signal C206: std_logic;
signal S206: std_logic;
signal C207: std_logic;
signal S207: std_logic;
signal C208: std_logic;
signal S208: std_logic;
signal C209: std_logic;
signal S209: std_logic;

begin

process(A,B)
begin

P0_0 <= A(0) AND B(0);
P1_0 <= A(1) AND B(0);
P2_0 <= A(2) AND B(0);
P3_0 <= A(3) AND B(0);
P4_0 <= A(4) AND B(0);
P5_0 <= A(5) AND B(0);
P6_0 <= A(6) AND B(0);
P7_0 <= A(7) AND B(0);
P8_0 <= A(8) AND B(0);
P9_0 <= A(9) AND B(0);
P10_0 <= A(10) AND B(0);
P11_0 <= A(11) AND B(0);
P12_0 <= A(12) AND B(0);
P13_0 <= A(13) AND B(0);
P14_0 <= A(14) AND B(0);
P0_1 <= A(0) AND B(1);
P1_1 <= A(1) AND B(1);
P2_1 <= A(2) AND B(1);
P3_1 <= A(3) AND B(1);
P4_1 <= A(4) AND B(1);
P5_1 <= A(5) AND B(1);
P6_1 <= A(6) AND B(1);
P7_1 <= A(7) AND B(1);
P8_1 <= A(8) AND B(1);
P9_1 <= A(9) AND B(1);
P10_1 <= A(10) AND B(1);
P11_1 <= A(11) AND B(1);
P12_1 <= A(12) AND B(1);
P13_1 <= A(13) AND B(1);
P14_1 <= A(14) AND B(1);
P0_2 <= A(0) AND B(2);
P1_2 <= A(1) AND B(2);
P2_2 <= A(2) AND B(2);
P3_2 <= A(3) AND B(2);
P4_2 <= A(4) AND B(2);
P5_2 <= A(5) AND B(2);
P6_2 <= A(6) AND B(2);
P7_2 <= A(7) AND B(2);
P8_2 <= A(8) AND B(2);
P9_2 <= A(9) AND B(2);
P10_2 <= A(10) AND B(2);
P11_2 <= A(11) AND B(2);
P12_2 <= A(12) AND B(2);
P13_2 <= A(13) AND B(2);
P14_2 <= A(14) AND B(2);
P0_3 <= A(0) AND B(3);
P1_3 <= A(1) AND B(3);
P2_3 <= A(2) AND B(3);
P3_3 <= A(3) AND B(3);
P4_3 <= A(4) AND B(3);
P5_3 <= A(5) AND B(3);
P6_3 <= A(6) AND B(3);
P7_3 <= A(7) AND B(3);
P8_3 <= A(8) AND B(3);
P9_3 <= A(9) AND B(3);
P10_3 <= A(10) AND B(3);
P11_3 <= A(11) AND B(3);
P12_3 <= A(12) AND B(3);
P13_3 <= A(13) AND B(3);
P14_3 <= A(14) AND B(3);
P0_4 <= A(0) AND B(4);
P1_4 <= A(1) AND B(4);
P2_4 <= A(2) AND B(4);
P3_4 <= A(3) AND B(4);
P4_4 <= A(4) AND B(4);
P5_4 <= A(5) AND B(4);
P6_4 <= A(6) AND B(4);
P7_4 <= A(7) AND B(4);
P8_4 <= A(8) AND B(4);
P9_4 <= A(9) AND B(4);
P10_4 <= A(10) AND B(4);
P11_4 <= A(11) AND B(4);
P12_4 <= A(12) AND B(4);
P13_4 <= A(13) AND B(4);
P14_4 <= A(14) AND B(4);
P0_5 <= A(0) AND B(5);
P1_5 <= A(1) AND B(5);
P2_5 <= A(2) AND B(5);
P3_5 <= A(3) AND B(5);
P4_5 <= A(4) AND B(5);
P5_5 <= A(5) AND B(5);
P6_5 <= A(6) AND B(5);
P7_5 <= A(7) AND B(5);
P8_5 <= A(8) AND B(5);
P9_5 <= A(9) AND B(5);
P10_5 <= A(10) AND B(5);
P11_5 <= A(11) AND B(5);
P12_5 <= A(12) AND B(5);
P13_5 <= A(13) AND B(5);
P14_5 <= A(14) AND B(5);
P0_6 <= A(0) AND B(6);
P1_6 <= A(1) AND B(6);
P2_6 <= A(2) AND B(6);
P3_6 <= A(3) AND B(6);
P4_6 <= A(4) AND B(6);
P5_6 <= A(5) AND B(6);
P6_6 <= A(6) AND B(6);
P7_6 <= A(7) AND B(6);
P8_6 <= A(8) AND B(6);
P9_6 <= A(9) AND B(6);
P10_6 <= A(10) AND B(6);
P11_6 <= A(11) AND B(6);
P12_6 <= A(12) AND B(6);
P13_6 <= A(13) AND B(6);
P14_6 <= A(14) AND B(6);
P0_7 <= A(0) AND B(7);
P1_7 <= A(1) AND B(7);
P2_7 <= A(2) AND B(7);
P3_7 <= A(3) AND B(7);
P4_7 <= A(4) AND B(7);
P5_7 <= A(5) AND B(7);
P6_7 <= A(6) AND B(7);
P7_7 <= A(7) AND B(7);
P8_7 <= A(8) AND B(7);
P9_7 <= A(9) AND B(7);
P10_7 <= A(10) AND B(7);
P11_7 <= A(11) AND B(7);
P12_7 <= A(12) AND B(7);
P13_7 <= A(13) AND B(7);
P14_7 <= A(14) AND B(7);
P0_8 <= A(0) AND B(8);
P1_8 <= A(1) AND B(8);
P2_8 <= A(2) AND B(8);
P3_8 <= A(3) AND B(8);
P4_8 <= A(4) AND B(8);
P5_8 <= A(5) AND B(8);
P6_8 <= A(6) AND B(8);
P7_8 <= A(7) AND B(8);
P8_8 <= A(8) AND B(8);
P9_8 <= A(9) AND B(8);
P10_8 <= A(10) AND B(8);
P11_8 <= A(11) AND B(8);
P12_8 <= A(12) AND B(8);
P13_8 <= A(13) AND B(8);
P14_8 <= A(14) AND B(8);
P0_9 <= A(0) AND B(9);
P1_9 <= A(1) AND B(9);
P2_9 <= A(2) AND B(9);
P3_9 <= A(3) AND B(9);
P4_9 <= A(4) AND B(9);
P5_9 <= A(5) AND B(9);
P6_9 <= A(6) AND B(9);
P7_9 <= A(7) AND B(9);
P8_9 <= A(8) AND B(9);
P9_9 <= A(9) AND B(9);
P10_9 <= A(10) AND B(9);
P11_9 <= A(11) AND B(9);
P12_9 <= A(12) AND B(9);
P13_9 <= A(13) AND B(9);
P14_9 <= A(14) AND B(9);
P0_10 <= A(0) AND B(10);
P1_10 <= A(1) AND B(10);
P2_10 <= A(2) AND B(10);
P3_10 <= A(3) AND B(10);
P4_10 <= A(4) AND B(10);
P5_10 <= A(5) AND B(10);
P6_10 <= A(6) AND B(10);
P7_10 <= A(7) AND B(10);
P8_10 <= A(8) AND B(10);
P9_10 <= A(9) AND B(10);
P10_10 <= A(10) AND B(10);
P11_10 <= A(11) AND B(10);
P12_10 <= A(12) AND B(10);
P13_10 <= A(13) AND B(10);
P14_10 <= A(14) AND B(10);
P0_11 <= A(0) AND B(11);
P1_11 <= A(1) AND B(11);
P2_11 <= A(2) AND B(11);
P3_11 <= A(3) AND B(11);
P4_11 <= A(4) AND B(11);
P5_11 <= A(5) AND B(11);
P6_11 <= A(6) AND B(11);
P7_11 <= A(7) AND B(11);
P8_11 <= A(8) AND B(11);
P9_11 <= A(9) AND B(11);
P10_11 <= A(10) AND B(11);
P11_11 <= A(11) AND B(11);
P12_11 <= A(12) AND B(11);
P13_11 <= A(13) AND B(11);
P14_11 <= A(14) AND B(11);
P0_12 <= A(0) AND B(12);
P1_12 <= A(1) AND B(12);
P2_12 <= A(2) AND B(12);
P3_12 <= A(3) AND B(12);
P4_12 <= A(4) AND B(12);
P5_12 <= A(5) AND B(12);
P6_12 <= A(6) AND B(12);
P7_12 <= A(7) AND B(12);
P8_12 <= A(8) AND B(12);
P9_12 <= A(9) AND B(12);
P10_12 <= A(10) AND B(12);
P11_12 <= A(11) AND B(12);
P12_12 <= A(12) AND B(12);
P13_12 <= A(13) AND B(12);
P14_12 <= A(14) AND B(12);
P0_13 <= A(0) AND B(13);
P1_13 <= A(1) AND B(13);
P2_13 <= A(2) AND B(13);
P3_13 <= A(3) AND B(13);
P4_13 <= A(4) AND B(13);
P5_13 <= A(5) AND B(13);
P6_13 <= A(6) AND B(13);
P7_13 <= A(7) AND B(13);
P8_13 <= A(8) AND B(13);
P9_13 <= A(9) AND B(13);
P10_13 <= A(10) AND B(13);
P11_13 <= A(11) AND B(13);
P12_13 <= A(12) AND B(13);
P13_13 <= A(13) AND B(13);
P14_13 <= A(14) AND B(13);
P0_14 <= A(0) AND B(14);
P1_14 <= A(1) AND B(14);
P2_14 <= A(2) AND B(14);
P3_14 <= A(3) AND B(14);
P4_14 <= A(4) AND B(14);
P5_14 <= A(5) AND B(14);
P6_14 <= A(6) AND B(14);
P7_14 <= A(7) AND B(14);
P8_14 <= A(8) AND B(14);
P9_14 <= A(9) AND B(14);
P10_14 <= A(10) AND B(14);
P11_14 <= A(11) AND B(14);
P12_14 <= A(12) AND B(14);
P13_14 <= A(13) AND B(14);
P14_14 <= A(14) AND B(14);

if ((A(15)='1' and B(15)='1') or (A(15)='0' and B(15)='0')) then
O(29) <= '0';
elsif ((A(15)='1' and B(15)='0') or (A(15)='0' and B(15)='1')) then
O(29) <= '1';
end if;

end process;

O(0) <= P0_0; 

FA1: Full_Adder port map(P1_0, P0_1, '0', S0, C0);

O(1) <= S0;

FA2: Full_Adder port map(P2_0, P1_1, P0_2, S1, C1);
FA3: Full_Adder port map(S1, C0, '0', S2, C2);

O(2) <= S2;

FA4: Full_Adder port map(P3_0, P2_1, P1_2, S3, C3);
FA5: Full_Adder port map(S3, P0_3, C2, S4, C4);
FA6: Full_Adder port map(S4, C1, '0', S5, C5);

O(3) <= S5;

FA7: Full_Adder port map(P4_0, P3_1, P2_2, S6, C6);
FA8: Full_Adder port map(S6, P1_3, P0_4, S7, C7);
FA9: Full_Adder port map(S7, C3, C4, S8, C8);
FA10: Full_Adder port map(S8, C5, '0', S9, C9);

O(4) <= S9;

FA11: Full_Adder port map(P5_0, P4_1, P3_2, S10, C10);
FA12: Full_Adder port map(P2_3, P1_4, P0_5, S11, C11);
FA13: Full_Adder port map(S10, S11, C6, S12, C12);
FA14: Full_Adder port map(S12, C7, C8, S13, C13);
FA15: Full_Adder port map(S13, C9, '0', S14, C14);

O(5) <= S14;

FA16: Full_Adder port map(P6_0, P5_1, P4_2, S15, C15);
FA17: Full_Adder port map(S15, P3_3, P2_4, S16, C16);
FA18: Full_Adder port map(S16, P1_5, P0_6, S17, C17);
FA19: Full_Adder port map(S17, C10, C11, S18, C18);
FA20: Full_Adder port map(S18, C12, C13, S19, C19);
FA21: Full_Adder port map(S19, C14, '0', S20, C20);

O(6) <= S20;

FA22: Full_Adder port map(P7_0, P6_1, P5_2, S21, C21);
FA23: Full_Adder port map(S21, P4_3, P3_4, S22, C22);
FA24: Full_Adder port map(S22, P2_5, P1_6, S23, C23);
FA25: Full_Adder port map(S23, P0_7, C15, S24, C24);
FA26: Full_Adder port map(S24, C16, C17, S25, C25);
FA27: Full_Adder port map(S25, C18, C19, S26, C26);
FA28: Full_Adder port map(S26, C20, '0', S27, C27);

O(7) <= S27;

FA29: Full_Adder port map(P8_0, P7_1, P6_2, S28, C28);
FA30: Full_Adder port map(S28, P5_3, P4_4, S29, C29);
FA31: Full_Adder port map(S29, P3_5, P2_6, S30, C30);
FA32: Full_Adder port map(S30, P1_7, P0_8, S31, C31);
FA33: Full_Adder port map(S31, C21, C22, S32, C32);
FA34: Full_Adder port map(S32, C23, C24, S33, C33);
FA35: Full_Adder port map(S33, C25, C26, S34, C34);
FA36: Full_Adder port map(S34, C27, '0', S35, C35);

O(8) <= S35;

FA37: Full_Adder port map(P9_0, P8_1, P7_2, S36, C36);
FA38: Full_Adder port map(S36, P6_3, P5_4, S37, C37);
FA39: Full_Adder port map(S37, P4_5, P3_6, S38, C38);
FA40: Full_Adder port map(S38, P2_7, P1_8, S39, C39);
FA41: Full_Adder port map(S39, P0_9, C28, S40, C40);
FA42: Full_Adder port map(S40, C29, C30, S41, C41);
FA43: Full_Adder port map(S41, C31, C32, S42, C42);
FA44: Full_Adder port map(S42, C33, C34, S43, C43);
FA45: Full_Adder port map(S43, C35, '0', S44, C44);

O(9) <= S44;

FA46: Full_Adder port map(P10_0, P9_1, P8_2, S45, C45);
FA47: Full_Adder port map(S45, P7_3, P6_4, S46, C46);
FA48: Full_Adder port map(S46, P5_5, P4_6, S47, C47);
FA49: Full_Adder port map(S47, P3_7, P2_8, S48, C48);
FA50: Full_Adder port map(S48, P1_9, P0_10, S49, C49);
FA51: Full_Adder port map(S49, C36, C37, S50, C50);
FA52: Full_Adder port map(S50, C38, C39, S51, C51);
FA53: Full_Adder port map(S51, C40, C41, S52, C52);
FA54: Full_Adder port map(S52, C42, C43, S53, C53);
FA55: Full_Adder port map(S53, C44, '0', S54, C54);

O(10) <= S54;

FA56: Full_Adder port map(P11_0, P10_1, P9_2, S55, C55);
FA57: Full_Adder port map(S55, P8_3, P7_4, S56, C56);
FA58: Full_Adder port map(S56, P6_5, P5_6, S57, C57);
FA59: Full_Adder port map(S57, P4_7, P3_8, S58, C58);
FA60: Full_Adder port map(S58, P2_9, P1_10, S59, C59);
FA61: Full_Adder port map(S59, P0_11, C45, S60, C60);
FA62: Full_Adder port map(S60, C46, C47, S61, C61);
FA63: Full_Adder port map(S61, C48, C49, S62, C62);
FA64: Full_Adder port map(S62, C50, C51, S63, C63);
FA65: Full_Adder port map(S63, C52, C53, S64, C64);
FA66: Full_Adder port map(S64, C54, '0', S65, C65);

O(11) <= S65;

FA67: Full_Adder port map(P12_0, P11_1, P10_2, S66, C66);
FA68: Full_Adder port map(S66, P9_3, P8_4, S67, C67);
FA69: Full_Adder port map(S67, P7_5, P6_6, S68, C68);
FA70: Full_Adder port map(S68, P5_7, P4_8, S69, C69);
FA71: Full_Adder port map(S69, P3_9, P2_10, S70, C70);
FA72: Full_Adder port map(S70, P1_11, P0_12, S71, C71);
FA73: Full_Adder port map(S71, C55, C56, S72, C72);
FA74: Full_Adder port map(S72, C57, C58, S73, C73);
FA75: Full_Adder port map(S73, C59, C60, S74, C74);
FA76: Full_Adder port map(S74, C61, C62, S75, C75);
FA77: Full_Adder port map(S75, C63, C64, S76, C76);
FA78: Full_Adder port map(S76, C65, '0', S77, C77);

O(12) <= S77;

FA79: Full_Adder port map(P13_0, P12_1, P11_2, S78, C78);
FA80: Full_Adder port map(S78, P10_3, P9_4, S79, C79);
FA81: Full_Adder port map(S79, P8_5, P7_6, S80, C80);
FA82: Full_Adder port map(S80, P6_7, P5_8, S81, C81);
FA83: Full_Adder port map(S81, P4_9, P3_10, S82, C82);
FA84: Full_Adder port map(S82, P2_11, P1_12, S83, C83);
FA85: Full_Adder port map(S83, P0_13, C66, S84, C84);
FA86: Full_Adder port map(S84, C67, C68, S85, C85);
FA87: Full_Adder port map(S85, C69, C70, S86, C86);
FA88: Full_Adder port map(S86, C71, C72, S87, C87);
FA89: Full_Adder port map(S87, C73, C74, S88, C88);
FA90: Full_Adder port map(S88, C75, C76, S89, C89);
FA91: Full_Adder port map(S89, C77, '0', S90, C90);

O(13) <= S90;

FA92: Full_Adder port map(P14_0, P13_1, P12_2, S91, C91);
FA93: Full_Adder port map(S91, P11_3, P10_4, S92, C92);
FA94: Full_Adder port map(S92, P9_5, P8_6, S93, C93);
FA95: Full_Adder port map(S93, P7_7, P6_8, S94, C94);
FA96: Full_Adder port map(S94, P5_9, P4_10, S95, C95);
FA97: Full_Adder port map(S95, P3_11, P2_12, S96, C96);
FA98: Full_Adder port map(S96, P1_13, P0_14, S97, C97);
FA99: Full_Adder port map(S97, C78, C79, S98, C98);
FA100: Full_Adder port map(S98, C80, C81, S99, C99);
FA101: Full_Adder port map(S99, C82, C83, S100, C100);
FA102: Full_Adder port map(S100, C84, C85, S101, C101);
FA103: Full_Adder port map(S101, C86, C87, S102, C102);
FA104: Full_Adder port map(S102, C88, C89, S103, C103);
FA105: Full_Adder port map(S103, C90, '0', S104, C104);

O(14) <= S104;

FA106: Full_Adder port map(P14_1, P13_2, P12_3, S105, C105);
FA107: Full_Adder port map(S105, P11_4, P10_5, S106, C106);
FA108: Full_Adder port map(S106, P9_6, P8_7, S107, C107);
FA109: Full_Adder port map(S107, P7_8, P6_9, S108, C108);
FA110: Full_Adder port map(S108, P5_10, P4_11, S109, C109);
FA111: Full_Adder port map(S109, P3_12, P2_13, S110, C110);
FA112: Full_Adder port map(S110, P1_14, C91, S111, C111);
FA113: Full_Adder port map(S111, C92, C93, S112, C112);
FA114: Full_Adder port map(S112, C94, C95, S113, C113);
FA115: Full_Adder port map(S113, C96, C97, S114, C114);
FA116: Full_Adder port map(S114, C98, C99, S115, C115);
FA117: Full_Adder port map(S115, C100, C101, S116, C116);
FA118: Full_Adder port map(S116, C102, C103, S117, C117);
FA119: Full_Adder port map(S117, C104, '0', S118, C118);

O(15) <= S118;

FA120: Full_Adder port map(P14_2, P13_3, P12_4, S119, C119);
FA121: Full_Adder port map(S119, P11_5, P10_6, S120, C120);
FA122: Full_Adder port map(S120, P9_7, P8_8, S121, C121);
FA123: Full_Adder port map(S121, P7_9, P6_10, S122, C122);
FA124: Full_Adder port map(S122, P5_11, P4_12, S123, C123);
FA125: Full_Adder port map(S123, P3_13, P2_14, S124, C124);
FA126: Full_Adder port map(S124, C105, C106, S125, C125);
FA127: Full_Adder port map(S125, C107, C108, S126, C126);
FA128: Full_Adder port map(S126, C109, C110, S127, C127);
FA129: Full_Adder port map(S127, C111, C112, S128, C128);
FA130: Full_Adder port map(S128, C113, C114, S129, C129);
FA131: Full_Adder port map(S129, C115, C116, S130, C130);
FA132: Full_Adder port map(S130, C117, C118, S131, C131);

O(16) <= S131;

FA133: Full_Adder port map(P14_3, P13_4, P12_5, S132, C132);
FA134: Full_Adder port map(S132, P11_6, P10_7, S133, C133);
FA135: Full_Adder port map(S133, P9_8, P8_9, S134, C134);
FA136: Full_Adder port map(S134, P7_10, P6_11, S135, C135);
FA137: Full_Adder port map(S135, P5_12, P4_13, S136, C136);
FA138: Full_Adder port map(S136, P3_14, C119, S137, C137);
FA139: Full_Adder port map(S137, C120, C121, S138, C138);
FA140: Full_Adder port map(S138, C122, C123, S139, C139);
FA141: Full_Adder port map(S139, C124, C125, S140, C140);
FA142: Full_Adder port map(S140, C126, C127, S141, C141);
FA143: Full_Adder port map(S141, C128, C129, S142, C142);
FA144: Full_Adder port map(S142, C130, C131, S143, C143);

O(17) <= S143;

FA145: Full_Adder port map(P14_4, P13_5, P12_6, S144, C144);
FA146: Full_Adder port map(S144, P11_7, P10_8, S145, C145);
FA147: Full_Adder port map(S145, P9_9, P8_10, S146, C146);
FA148: Full_Adder port map(S146, P7_11, P6_12, S147, C147);
FA149: Full_Adder port map(S147, P5_13, P4_14, S148, C148);
FA150: Full_Adder port map(S148, C132, C133, S149, C149);
FA151: Full_Adder port map(S149, C134, C135, S150, C150);
FA152: Full_Adder port map(S150, C136, C137, S151, C151);
FA153: Full_Adder port map(S151, C138, C139, S152, C152);
FA154: Full_Adder port map(S152, C140, C141, S153, C153);
FA155: Full_Adder port map(S153, C142, C143, S154, C154);

O(18) <= S154;

FA156: Full_Adder port map(P14_5, P13_6, P12_7, S155, C155);
FA157: Full_Adder port map(S155, P11_8, P10_9, S156, C156);
FA158: Full_Adder port map(S156, P9_10, P8_11, S157, C157);
FA159: Full_Adder port map(S157, P7_12, P6_13, S158, C158);
FA160: Full_Adder port map(S158, P5_14, C144, S159, C159);
FA161: Full_Adder port map(S159, C145, C146, S160, C160);
FA162: Full_Adder port map(S160, C147, C148, S161, C161);
FA163: Full_Adder port map(S161, C149, C150, S162, C162);
FA164: Full_Adder port map(S162, C151, C152, S163, C163);
FA165: Full_Adder port map(S163, C153, C154, S164, C164);

O(19) <= S164;

FA166: Full_Adder port map(P14_6, P13_7, P12_8, S165, C165);
FA167: Full_Adder port map(S165, P11_9, P10_10, S166, C166);
FA168: Full_Adder port map(S166, P9_11, P8_12, S167, C167);
FA169: Full_Adder port map(S167, P7_13, P6_14, S168, C168);
FA170: Full_Adder port map(S168, C155, C156, S169, C169);
FA171: Full_Adder port map(S169, C157, C158, S170, C170);
FA172: Full_Adder port map(S170, C159, C160, S171, C171);
FA173: Full_Adder port map(S171, C161, C162, S172, C172);
FA174: Full_Adder port map(S172, C163, C164, S173, C173);

O(20) <= S173;

FA175: Full_Adder port map(P14_7, P13_8, P12_9, S174, C174);
FA176: Full_Adder port map(S174, P11_10, P10_11, S175, C175);
FA177: Full_Adder port map(S175, P9_12, P8_13, S176, C176);
FA178: Full_Adder port map(S176, P7_14, C165, S177, C177);
FA179: Full_Adder port map(S177, C166, C167, S178, C178);
FA180: Full_Adder port map(S178, C168, C169, S179, C179);
FA181: Full_Adder port map(S179, C170, C171, S180, C180);
FA182: Full_Adder port map(S180, C172, C173, S181, C181);

O(21) <= S181;

FA183: Full_Adder port map(P14_8, P13_9, P12_10, S182, C182);
FA184: Full_Adder port map(S182, P11_11, P10_12, S183, C183);
FA185: Full_Adder port map(S183, P9_13, P8_14, S184, C184);
FA186: Full_Adder port map(S184, C174, C175, S185, C185);
FA187: Full_Adder port map(S185, C176, C177, S186, C186);
FA188: Full_Adder port map(S186, C178, C179, S187, C187);
FA189: Full_Adder port map(S187, C180, C181, S188, C188);

O(22) <= S188;

FA190: Full_Adder port map(P14_9, P13_10, P12_11, S189, C189);
FA191: Full_Adder port map(S189, P11_12, P10_13, S190, C190);
FA192: Full_Adder port map(S190, P9_14, C182, S191, C191);
FA193: Full_Adder port map(S191, C183, C184, S192, C192);
FA194: Full_Adder port map(S192, C185, C186, S193, C193);
FA195: Full_Adder port map(S193, C187, C188, S194, C194);

O(23) <= S194;

FA196: Full_Adder port map(P14_10, P13_11, P12_12, S195, C195);
FA197: Full_Adder port map(S195, P11_13, P10_14, S196, C196);
FA198: Full_Adder port map(S196, C189, C190, S197, C197);
FA199: Full_Adder port map(S197, C191, C192, S198, C198);
FA200: Full_Adder port map(S198, C193, C194, S199, C199);

O(24) <= S199;

FA201: Full_Adder port map(P14_11, P13_12, P12_13, S200, C200);
FA202: Full_Adder port map(S200, P11_14, C195, S201, C201);
FA203: Full_Adder port map(S201, C196, C197, S202, C202);
FA204: Full_Adder port map(S202, C198, C199, S203, C203);

O(25) <= S203;

FA205: Full_Adder port map(P14_12, P13_13, P12_14, S204, C204);
FA206: Full_Adder port map(S204, C200, C201, S205, C205);
FA207: Full_Adder port map(S205, C202, C203, S206, C206);

O(26) <= S206;

FA208: Full_Adder port map(P14_13, P13_14, C204, S207, C207);
FA209: Full_Adder port map(S207, C205, C206, S208, C208);

O(27) <= S208;

FA210: Full_Adder port map(P14_14, C207, C208, S209, C209);

O(28) <= S209;

end Behavioral;
